module main

import term.ui as tui

const (
	white = tui.Color{
		r: 240
		g: 240
		b: 240
	}
	blue = tui.Color{
		r: 100
		g: 220
		b: 220
	}
	red = tui.Color{
		r: 200
		g: 0
		b: 0
	}
	grey = tui.Color{
		r: 200
		g: 200
		b: 200
	}
	black = tui.Color{
		r: 10
		g: 10
		b: 10
	}
)
